package test_pkg;
  import uvm_pkg::*;

  `include "btb_seq_item.sv"
  `include "btb_sequencer.sv"
  `include "btb_driver.sv"
  `include "btb_monitor.sv"
  `include "btb_agent.sv"
  `include "btb_scoreboard.sv"
  `include "btb_env.sv"
  `include "btb_test.sv"
  `include "btb_generic_test.sv"

endpackage
